// AUTO CODE, don't edit!
//   
module __MOD_NAME__
    #(parameter BASE_ADDR=0
    input               rst,

    input     [__BUS_AWID__-1:0]  bif_addr,
    //__ ITR_FIELD:PORT DEF BEGIN(py:ctx['field']['attr']['acc']['type']=='intact' or ctx['field']['split_idx']==0)
    __SIG_DIR__ __SIG_WID_DEF__ __SIG_NAME__,
    //__ ITR_FIELD:PORT DEF END

    // dummy
    output              tie0

